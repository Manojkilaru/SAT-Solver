-- This testbench will result in an unsat condition.In this testbench we gave 1024 clauses. 
--The stress in this testbench is that we varied the first 10 variabels giving all the 2^10 possible clauses for these 10 variables 
--and assigning 0's to all the other variables from x11-64. This test case checks the 2^10 possible cases i.e., it runs in 2^10 clock cycles
--(In our system the sat became 0 at t = 30,855ns).


--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   23:32:12 04/06/2016
-- Design Name:   
-- Module Name:   C:/Users/chanukya/Desktop/Xilinx/SATSolver/Pirates_testbench1.vhd
-- Project Name:  SATSolver
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Input
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Pirates_testbench1 IS
END Pirates_testbench1;
 
ARCHITECTURE behavior OF Pirates_testbench1 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Input
    PORT(
         clock : IN  std_logic;
         reset : IN  std_logic;
         clause : IN  std_logic_vector(63 downto 0);
         load : IN  std_logic;
         SAT : INOUT  std_logic;
         output : INOUT  std_logic_vector(63 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clock : std_logic := '0';
   signal reset : std_logic := '0';
   signal clause : std_logic_vector(63 downto 0) := (others => '0');
   signal load : std_logic := '0';

	--BiDirs
   signal SAT : std_logic;
   signal output : std_logic_vector(63 downto 0);

   -- Clock period definitions
   constant clock_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Input PORT MAP (
          clock => clock,
          reset => reset,
          clause => clause,
          load => load,
          SAT => SAT,
          output => output
        );

   -- Clock process definitions
   clock_process :process
   begin
		clock <= '0';
		wait for clock_period/2;
		clock <= '1';
		wait for clock_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;
		reset <= '1';
		wait for 2*clock_period;
		reset <= '0';
			load<='1';
		clause<="0000000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1000111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0111000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1001111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0110000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1010111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0101000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1011111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0100000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1100111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0011000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1101111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0010000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1110111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0001000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111100111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000011000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111101111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000010000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111110111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000001000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111100000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000011000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111101000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000010000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111110000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000001000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="1111111111000000000000000000000000000000000000000000000000000000";
		wait for clock_period;
	load<='1';
		clause<="0000000000000000000000000000000000000000000000000000000000000000";
		wait for clock_period;

		load<='0';

      wait;
   end process;

END;
